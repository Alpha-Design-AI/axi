// TODO: Implement the axi_to_axi_lite module here
// See TASK.md and test/tb_axi_to_axi_lite.sv for requirements

module axi_to_axi_lite #(
    // Add your parameters here
) (
    // Add your ports here
);
    // Add your implementation here
endmodule
