// TODO: Implement the axi_modify_address module here
// See TASK.md and test/tb_axi_modify_address.sv for requirements

module axi_modify_address #(
    // Add your parameters here
) (
    // Add your ports here
);
    // Add your implementation here
endmodule
