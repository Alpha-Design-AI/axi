// TODO: Implement the axi_atop_filter module here
// See TASK.md and test/tb_axi_atop_filter.sv for requirements

module axi_atop_filter #(
    // Add your parameters here
) (
    // Add your ports here
);
    // Add your implementation here
endmodule
