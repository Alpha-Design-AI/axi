// TODO: Implement the axi_iw_converter module here
// See TASK.md and test/tb_axi_iw_converter.sv for requirements

module axi_iw_converter #(
    // Add your parameters here
) (
    // Add your ports here
);
    // Add your implementation here
endmodule
