// TODO: Implement the axi_lite_regs module here
// See TASK.md and test/tb_axi_lite_regs.sv for requirements

module axi_lite_regs #(
    // Add your parameters here
) (
    // Add your ports here
);
    // Add your implementation here
endmodule
