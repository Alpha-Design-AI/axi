// TODO: Implement the axi_sim_mem module here
// See TASK.md and test/tb_axi_sim_mem.sv for requirements

module axi_sim_mem #(
    // Add your parameters here
) (
    // Add your ports here
);
    // Add your implementation here
endmodule
