// TODO: Implement the axi_isolate module here
// See TASK.md and test/tb_axi_isolate.sv for requirements

module axi_isolate #(
    // Add your parameters here
) (
    // Add your ports here
);
    // Add your implementation here
endmodule
