// TODO: Implement the axi_lite_mailbox module here
// See TASK.md and test/tb_axi_lite_mailbox.sv for requirements

module axi_lite_mailbox #(
    // Add your parameters here
) (
    // Add your ports here
);
    // Add your implementation here
endmodule
