// TODO: Implement the axi_delayer module here
// See TASK.md and test/tb_axi_delayer.sv for requirements

module axi_delayer #(
    // Add your parameters here
) (
    // Add your ports here
);
    // Add your implementation here
endmodule
