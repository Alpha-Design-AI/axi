// TODO: Implement the axi_serializer module here
// See TASK.md and test/tb_axi_serializer.sv for requirements

module axi_serializer #(
    // Add your parameters here
) (
    // Add your ports here
);
    // Add your implementation here
endmodule
