// TODO: Implement the axi_lite_to_axi module here
// See TASK.md and test/tb_axi_lite_to_axi.sv for requirements

module axi_lite_to_axi #(
    // Add your parameters here
) (
    // Add your ports here
);
    // Add your implementation here
endmodule
