// TODO: Implement the axi_fifo module here
// See TASK.md and test/tb_axi_fifo.sv for requirements

module axi_fifo #(
    // Add your parameters here
) (
    // Add your ports here
);
    // Add your implementation here
endmodule
